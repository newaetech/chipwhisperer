/***********************************************************************
This file is part of the ChipWhisperer Project. See www.newae.com for more
details, or the codebase at http://www.chipwhisperer.com

Copyright (c) 2022, NewAE Technology Inc. All rights reserved.
Author: Jean-Pierre Thibault <jpthibault@newae.com>

  chipwhisperer is free software: you can redistribute it and/or modify
  it under the terms of the GNU General Public License as published by
  the Free Software Foundation, either version 3 of the License, or
  (at your option) any later version.

  chipwhisperer is distributed in the hope that it will be useful,
  but WITHOUT ANY WARRANTY; without even the implied warranty of
  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
  GNU Lesser General Public License for more details.

  You should have received a copy of the GNU General Public License
  along with chipwhisperer.  If not, see <http://www.gnu.org/licenses/>.
*************************************************************************/

//////////////////////////////////////////////////////////////////////////////////
// General Top-Level Module for iCEUP5K Target. 
// Adapted from CW308T_S6LX9_SS.v.
//
//////////////////////////////////////////////////////////////////////////////////


`timescale 1 ns / 1ps
`default_nettype none

module iCE40UP5K_SS_example (
    input  wire cw_clk,         // 45A_G1 pin, header B
    input  wire ice_clk,
    input  wire clk_sel,        // 37A pin, SW2
    input  wire clk_alive_en,   // 36B pin, SW2
    output wire TxD,            // 42B pin, header B
    input  wire RxD,            // 43A pin, header B
    output wire IO4,            // 38B pin, header B
    output wire led_green,
    output wire led_blue,
    output wire led_red
);

    wire LED_rx;
    wire LED_go;

    assign led_green = ~(LED_rx & ~LED_go);
    assign led_red = ~(LED_go & ~LED_rx);
    assign led_blue = clk_alive_en? ~count[23] : 1'b1;

    reg [23:0] count;
    always @(posedge clk) count <= count + 1;

    wire [127:0] enc_input;     // Input to encryption algorithm (normally PT)
    wire [127:0] enc_output;    // Output from encryption algorithm (normally CT)
    wire [127:0] enc_key;       // Encryption key to use
    wire load_input;            // One-clock cycle flag to indicate data in enc_input is valid
    wire load_key;              // One-cycle flag to indicate data in enc_input is valid
    wire enc_go;                // One-cycle flag to indicate we should run an encryption
    wire enc_output_ready;      // One-cycle flag generated by encryption core indicating data out is valid

    wire clk = clk_sel? ice_clk : cw_clk;

    SimpleSerial SSCore(
        .clk            (clk), 
        .TxD            (TxD), 
        .RxD            (RxD), 
        .LED_rx         (LED_rx), 
        .LED_go         (LED_go),
        .pt             (enc_input), 
        .key            (enc_key), 
        .load_key       (load_key), 
        .load_pt        (load_input),
        .do_enc         (enc_go), 
        .ct             (enc_output), 
        .ct_ready       (enc_output_ready)
    );

    wire enc_busy;
    assign IO4 = enc_busy;

    aes_core AESGoogleVault(
        .clk        (clk),
        .load_i     (enc_go),
        .key_i      ({enc_key, 128'h0}),
        .data_i     (enc_input),
        .size_i     (2'd0),
        .dec_i      (1'b0),
        .data_o     (enc_output),
        .busy_o     (enc_busy)
    );

    //Generate single-clock cycle pulse when enc_busy falls
    reg enc_done_flag;
    reg enc_busy_delayed;

    always @(posedge clk) begin
        enc_busy_delayed <= enc_busy;
        enc_done_flag <= ~enc_busy & enc_busy_delayed;
    end

    assign enc_output_ready = enc_done_flag;

endmodule

`default_nettype wire

